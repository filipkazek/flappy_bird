
package vga_pkg;

  
    localparam HOR_PIXELS = 1024;
    localparam VER_PIXELS = 768;
    localparam HOR_TOTAL_TIME = 1344;
    localparam HOR_BLANK_TIME = 320;
    localparam HOR_SYNC_START = 1048;
    localparam HOR_SYNC_TIME = 136;
    localparam VER_TOTAL_TIME = 806;
    localparam VER_BLANK_TIME = 38;
    localparam VER_SYNC_START = 771;
    localparam VER_SYNC_TIME = 6;




endpackage
